`timescale 1ns/10ps
module test;

endmodule
